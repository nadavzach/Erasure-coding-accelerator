

module module_tb_wrapper#(

   //------------------------------------------
   //--- Interface Parameters:
   //------------------------------------------
   

   //------------------------------------------
   //---testbench Parameters:
   //------------------------------------------

   parameter CLK_CYC = 10

   
   );

  

    
    //General
    logic          clk;
    logic          rst_n;

    //Internal signals
    logic start;
    logic finish;
    //logics:
    //******************************************
    //
    //******************************************

  
   
  
   //******************************************
   //  output for TB and debugging
   //******************************************
  


   
 

 //#################################################            
// ================================================
// ~~~~~~~~~~ Instantiations ~~~~~~~~~~
// ================================================
//#################################################




                       
//******************************************
// Instantiation - "module name"
//******************************************
//input dly assignment 
//******************************************
assign #IF_DLY <signal name>_dly = <signal name>;
   
    

// ================================================
// ~~~~~~~~~~ test bench logic ~~~~~~~~~~
// ================================================

//Init
initial
begin
    clk		    	 <= 1'b0;
    rst_n            <= 1'b0;
    #(3*CLK_CYCLE) 
    
    rst_n <= 1'b1;
    

end

//-----------------------------------
//Clocks
//-----------------------------------

always
begin
    #(CLK_CYCLE/2) clk <= ~clk;
end

//-----------------------------------
//Reseting logics
//-----------------------------------

always @(posedge clk or negedge rst_n)
begin
    if(~rst_n)
    begin
    <signal name>       <=      1'b0;
   
    end
    else
	start                                <= 1'b1;
end



// ================================================
// ~~~~~~~~~~ test bench flow ~~~~~~~~~~
// ================================================



always @(finish)
begin
    if (finish)
        $finish;
end

 endmodule

 
